library verilog;
use verilog.vl_types.all;
entity test1_vlg_vec_tst is
end test1_vlg_vec_tst;
