library verilog;
use verilog.vl_types.all;
entity flow_led_vlg_vec_tst is
end flow_led_vlg_vec_tst;
