library verilog;
use verilog.vl_types.all;
entity flow_LED_vlg_vec_tst is
end flow_LED_vlg_vec_tst;
